LPM_COUNTER_VARIANT_inst : LPM_COUNTER_VARIANT PORT MAP (
		clk_en	 => clk_en_sig,
		clock	 => clock_sig,
		sclr	 => sclr_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
